library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;

entity ROM_176x4 is
  port (Clock : in std_logic;
  		CS_L : in std_logic;
        R_W  : in std_logic;
        Addr   : in std_logic_vector(7 downto 0);
        Data  : out std_logic_vector(3 downto 0));
end ROM_176x4;

architecture ROM_176x4_Arch of ROM_176x4 is
  type rom_type is array (0 to 175)
        of std_logic_vector (3 downto 0);
  signal ROM : rom_type;
  signal Read_Enable : std_logic;
begin

ROM(0) <= X"5";
ROM(1) <= X"0";
ROM(2) <= X"B";
ROM(3) <= X"3";
ROM(4) <= X"6";
ROM(5) <= X"7";
ROM(6) <= X"0";
ROM(7) <= X"D";
ROM(8) <= X"0";
ROM(9) <= X"B";
ROM(10) <= X"F";
ROM(11) <= X"0";
ROM(12) <= X"B";
ROM(13) <= X"4";
ROM(14) <= X"2";
ROM(15) <= X"6";
ROM(16) <= X"1";
ROM(17) <= X"D";
ROM(18) <= X"0";
ROM(19) <= X"B";
ROM(20) <= X"5";
ROM(21) <= X"0";
ROM(22) <= X"B";
ROM(23) <= X"1";
ROM(24) <= X"6";
ROM(25) <= X"F";
ROM(26) <= X"0";
ROM(27) <= X"B";
ROM(28) <= X"B";
ROM(29) <= X"2";
ROM(30) <= X"2";
ROM(31) <= X"9";
ROM(32) <= X"A";
ROM(33) <= X"0";
ROM(34) <= X"4";
ROM(35) <= X"2";
ROM(36) <= X"6";
ROM(37) <= X"1";
ROM(38) <= X"4";
ROM(39) <= X"2";
ROM(40) <= X"D";
ROM(41) <= X"0";
ROM(42) <= X"B";
ROM(43) <= X"5";
ROM(44) <= X"0";
ROM(45) <= X"B";
ROM(46) <= X"3";
ROM(47) <= X"6";
ROM(48) <= X"F";
ROM(49) <= X"0";
ROM(50) <= X"B";
ROM(51) <= X"7";
ROM(52) <= X"0";
ROM(53) <= X"4";
ROM(54) <= X"2";
ROM(55) <= X"F";
ROM(56) <= X"1";
ROM(57) <= X"B";
ROM(58) <= X"6";
ROM(59) <= X"7";
ROM(60) <= X"A";
ROM(61) <= X"6";
ROM(62) <= X"5";
ROM(63) <= X"6";
ROM(64) <= X"A";
ROM(65) <= X"4";
ROM(66) <= X"1";
ROM(67) <= X"D";
ROM(68) <= X"1";
ROM(69) <= X"B";
ROM(70) <= X"5";
ROM(71) <= X"0";
ROM(72) <= X"B";
ROM(73) <= X"3";
ROM(74) <= X"6";
ROM(75) <= X"F";
ROM(76) <= X"1";
ROM(77) <= X"B";
ROM(78) <= X"7";
ROM(79) <= X"0";
ROM(80) <= X"D";
ROM(81) <= X"0";
ROM(82) <= X"B";
ROM(83) <= X"9";
ROM(84) <= X"A";
ROM(85) <= X"0";
ROM(86) <= X"4";
ROM(87) <= X"1";
ROM(88) <= X"7";
ROM(89) <= X"0";
ROM(90) <= X"D";
ROM(91) <= X"1";
ROM(92) <= X"B";
ROM(93) <= X"D";
ROM(94) <= X"0";
ROM(95) <= X"B";
ROM(96) <= X"9";
ROM(97) <= X"A";
ROM(98) <= X"0";
ROM(99) <= X"F";
ROM(100) <= X"0";
ROM(101) <= X"B";
ROM(102) <= X"A";
ROM(103) <= X"A";
ROM(104) <= X"7";
ROM(105) <= X"6";
ROM(106) <= X"F";
ROM(107) <= X"4";
ROM(108) <= X"2";
ROM(109) <= X"D";
ROM(110) <= X"0";
ROM(111) <= X"B";
ROM(112) <= X"5";
ROM(113) <= X"0";
ROM(114) <= X"6";
ROM(115) <= X"8";
ROM(116) <= X"B";
ROM(117) <= X"A";
ROM(118) <= X"0";
ROM(119) <= X"9";
ROM(120) <= X"3";
ROM(121) <= X"6";
ROM(122) <= X"F";
ROM(123) <= X"1";
ROM(124) <= X"B";
ROM(125) <= X"A";
ROM(126) <= X"C";
ROM(127) <= X"8";
ROM(128) <= X"6";
ROM(129) <= X"F";
ROM(130) <= X"4";
ROM(131) <= X"1";
ROM(132) <= X"D";
ROM(133) <= X"1";
ROM(134) <= X"B";
ROM(135) <= X"7";
ROM(136) <= X"9";
ROM(137) <= X"9";
ROM(138) <= X"B";
ROM(139) <= X"6";
ROM(140) <= X"7";
ROM(141) <= X"9";
ROM(142) <= X"4";
ROM(143) <= X"1";
ROM(144) <= X"D";
ROM(145) <= X"1";
ROM(146) <= X"B";
ROM(147) <= X"7";
ROM(148) <= X"9";
ROM(149) <= X"9";
ROM(150) <= X"B";
ROM(151) <= X"6";
ROM(152) <= X"0";
ROM(153) <= X"0";
ROM(154) <= X"0";
ROM(155) <= X"0";
ROM(156) <= X"0";
ROM(157) <= X"0";
ROM(158) <= X"0";
ROM(159) <= X"0";
ROM(160) <= X"0";
ROM(161) <= X"0";
ROM(162) <= X"0";
ROM(163) <= X"0";
ROM(164) <= X"0";
ROM(165) <= X"0";
ROM(166) <= X"0";
ROM(167) <= X"0";
ROM(168) <= X"0";
ROM(169) <= X"0";
ROM(170) <= X"0";
ROM(171) <= X"0";
ROM(172) <= X"0";
ROM(173) <= X"0";
ROM(174) <= X"0";
ROM(175) <= X"0";
	Read_Enable <=  '0' when(CS_L='0' and R_W = '1') else '1';

	process (Clock)
	begin
		if(Clock='0') then
			if(Read_Enable = '0') then
			  Data  <= ROM(conv_integer(Addr));
		  	else
			  Data <= "ZZZZ";
	      	end if;
		else Data <= "ZZZZ";
		end if;

	end process;

	end ROM_176x4_Arch;
